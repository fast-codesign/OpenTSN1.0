/*========================================================================================================*\
          Filename : gc.v,gate control
            Author : peng jintao
       Description : Judge whether four queues(Q0��Q1��Q2��Q3) can be scheduled; transmit result to TS module.
	     Called by : 
  Revision History : 5/16/2019 Revision 1.0  peng jintao
                     mm/dd/yy
           Company : 662
============================================================================================================
          Comments :
\*========================================================================================================*/
`timescale 1ns/1ps

module gc#(
    parameter    PLATFORM = "xilinx"
)(
//clk & rst
input	wire			clk,
input	wire			rst_n,

//receive from MB
input	wire     [3:0]  in_gc_md_outport,
input	wire     [3:0]  in_gc_fifo_empty,     
input	wire     [6:0]  in_gc_pkt_len,

//receive from LCM
input	wire            in_gc_time_slot_flag,
input	wire     [31:0] in_gc_rate_limit,       //100*8ns(per clock)*(rate(bps)/8)*(10^-9)= rate*(10^-7)��add number of token per 800ns(100 clocks); the minimum committed information rate 10Mbps is allowed.

//receive from EBM
input	wire            in_gc_pkt_valid,

//receive from UDO
input	wire      [7:0]  pktout_usedw_0,
input	wire      [7:0]  pktout_usedw_1,

//transmit to TS
output	reg      [3:0]  out_gc_schedule_valid,
//receive from TS
input	wire            in_gc_q2_rden

);

//token bucken parameter
localparam TB_size = 12'h7FF;   //committed burst size is 2047 Byte.
reg  [11:0] RT;        //remaining tokens
reg  [11:0] CT;        //consume tokens,1Byte consumes 1 token.
reg  [6:0]  TB_cnt;    //timer of token bucken

wire [11:0] pkt_len;
assign pkt_len = {5'b0,in_gc_pkt_len}<<4;

//************************************************************
//                   Consume tokens
//************************************************************
always@(posedge clk or negedge rst_n) begin
    if(rst_n == 1'b0) begin
        CT <= 12'd0;		
    end
    else begin
		if(in_gc_q2_rden == 1'b1)begin
		    CT <= pkt_len;
		end
		else begin
		    CT <= 12'd0;
		end
    end
end

//************************************************************
//                    Count token
//************************************************************
always@(negedge clk or posedge rst_n) begin
    if(rst_n == 1'b0) begin
        RT <= 12'd0;
		TB_cnt <= 7'd0;
    end
    else begin
	    if(TB_cnt >= 7'd99)begin
		    TB_cnt <= 7'd0;
			if(RT + in_gc_rate_limit[11:0] - CT <= TB_size)begin
			    RT <= RT + in_gc_rate_limit[11:0] - CT;
			end
			else begin
			    RT <= TB_size;
			end
		end
		else begin
		    TB_cnt <= TB_cnt + 7'd1;
			RT <= RT - CT;
		end
    end
end

//************************************************************
//        Judge whether four queues can be scheduled
//************************************************************
reg [1:0] state;
reg       init_flag;   
localparam IDLE_S = 2'd0,
           JUDGE_QUEUE_S = 2'd1;
always@(posedge clk or negedge rst_n) begin
    if(rst_n == 1'b0) begin
        out_gc_schedule_valid <= 4'b0;
		init_flag <= 1'b1;
		state <= IDLE_S;
    end
    else begin
	    case(state)
            IDLE_S:begin
			    if(init_flag || in_gc_pkt_valid)begin
				    state <= JUDGE_QUEUE_S;    
				end
				else begin
				    state <= IDLE_S; 
				end
			end
            JUDGE_QUEUE_S:begin
			    if(|out_gc_schedule_valid[3:0])begin
				    out_gc_schedule_valid <= 4'b0;
					init_flag <= 1'b0;
					state <= IDLE_S;
                end					
                else begin
				    state <= JUDGE_QUEUE_S;
				    if(in_gc_time_slot_flag && (!in_gc_fifo_empty[0]) && ((!in_gc_md_outport[0] && (pktout_usedw_0 <= 20)) || (in_gc_md_outport[0] && (pktout_usedw_1 <= 20))))begin    //Judge whether Q0 queue can be scheduled
		                out_gc_schedule_valid[0] <= 1'b1;					
                    end
		            else begin
		                out_gc_schedule_valid[0] <= 1'b0;
		            end
					
				    if(!in_gc_time_slot_flag && (!in_gc_fifo_empty[1]) && ((!in_gc_md_outport[1] && (pktout_usedw_0 <= 20)) || (in_gc_md_outport[1] && (pktout_usedw_1 <= 20))))begin   //Judge whether Q1 queue can be scheduled
		                out_gc_schedule_valid[1] <= 1'b1;
                    end
		            else begin
		                out_gc_schedule_valid[1] <= 1'b0;
					end
					
					if((RT >= pkt_len) && (!in_gc_fifo_empty[2]) && ((!in_gc_md_outport[2] && (pktout_usedw_0 <= 20)) || (in_gc_md_outport[2] && (pktout_usedw_1 <= 20))))begin        //Judge whether Q2 queue can be scheduled
		                out_gc_schedule_valid[2] <= 1'b1;  					
                    end
		            else begin
		                out_gc_schedule_valid[2] <= 1'b0;
		            end
					
					if((!in_gc_fifo_empty[3]) && ((!in_gc_md_outport[3] && (pktout_usedw_0 <= 20)) || (in_gc_md_outport[3] && (pktout_usedw_1 <= 20))))begin                          //Judge whether Q3 queue can be scheduled
		                out_gc_schedule_valid[3] <= 1'b1;			
                    end
		            else begin
		                out_gc_schedule_valid[3] <= 1'b0;
		            end
				end
		    end
	    endcase
    end     
end        

endmodule